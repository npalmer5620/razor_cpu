`timescale 1ns / 1ps
// Nicholas Palmer | March 12, 2023

module control_v2(

    );
endmodule
